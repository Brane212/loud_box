module shout_1(
input clk_in,
output pll_step, shout_out);










endmodule